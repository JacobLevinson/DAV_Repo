module Lab_7(LEDs);
output [7:0] LEDs;

endmodule